LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

-- Gerador de pulso que, por padrão, gera um pequeno pulso à frequência de 2Hz a partir de um clock de entrada de 50MHz.

ENTITY PulseGenerator IS
    GENERIC (MAX : POSITIVE := 25_000_000);
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        pulse : OUT STD_LOGIC);
END PulseGenerator;

ARCHITECTURE Behavioral OF PulseGenerator IS
    SIGNAL s_cnt : NATURAL RANGE 0 TO MAX - 1;
BEGIN
    PROCESS (clock)
    BEGIN
        IF (rising_edge(clock)) THEN
            pulse <= '0';
            IF (reset = '1') THEN
                s_cnt <= 0;
            ELSE
                s_cnt <= s_cnt + 1;
                IF (s_cnt = MAX - 1) THEN
                    s_cnt <= 0;
                    pulse <= '1';
                END IF;
            END IF;
        END IF;
    END PROCESS;
END Behavioral;